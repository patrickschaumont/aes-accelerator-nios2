module tboxe3(input wire clk,
              input wire [7:0] a,
              output reg [31:0] q);

   always @(posedge clk)
     case (a)
	8'd0: q = 32'h6363a5c6;
	8'd1: q = 32'h7c7c84f8;
	8'd2: q = 32'h777799ee;
	8'd3: q = 32'h7b7b8df6;
	8'd4: q = 32'hf2f20dff;
	8'd5: q = 32'h6b6bbdd6;
	8'd6: q = 32'h6f6fb1de;
	8'd7: q = 32'hc5c55491;
	8'd8: q = 32'h30305060;
	8'd9: q = 32'h1010302;
	8'd10: q = 32'h6767a9ce;
	8'd11: q = 32'h2b2b7d56;
	8'd12: q = 32'hfefe19e7;
	8'd13: q = 32'hd7d762b5;
	8'd14: q = 32'hababe64d;
	8'd15: q = 32'h76769aec;
	8'd16: q = 32'hcaca458f;
	8'd17: q = 32'h82829d1f;
	8'd18: q = 32'hc9c94089;
	8'd19: q = 32'h7d7d87fa;
	8'd20: q = 32'hfafa15ef;
	8'd21: q = 32'h5959ebb2;
	8'd22: q = 32'h4747c98e;
	8'd23: q = 32'hf0f00bfb;
	8'd24: q = 32'hadadec41;
	8'd25: q = 32'hd4d467b3;
	8'd26: q = 32'ha2a2fd5f;
	8'd27: q = 32'hafafea45;
	8'd28: q = 32'h9c9cbf23;
	8'd29: q = 32'ha4a4f753;
	8'd30: q = 32'h727296e4;
	8'd31: q = 32'hc0c05b9b;
	8'd32: q = 32'hb7b7c275;
	8'd33: q = 32'hfdfd1ce1;
	8'd34: q = 32'h9393ae3d;
	8'd35: q = 32'h26266a4c;
	8'd36: q = 32'h36365a6c;
	8'd37: q = 32'h3f3f417e;
	8'd38: q = 32'hf7f702f5;
	8'd39: q = 32'hcccc4f83;
	8'd40: q = 32'h34345c68;
	8'd41: q = 32'ha5a5f451;
	8'd42: q = 32'he5e534d1;
	8'd43: q = 32'hf1f108f9;
	8'd44: q = 32'h717193e2;
	8'd45: q = 32'hd8d873ab;
	8'd46: q = 32'h31315362;
	8'd47: q = 32'h15153f2a;
	8'd48: q = 32'h4040c08;
	8'd49: q = 32'hc7c75295;
	8'd50: q = 32'h23236546;
	8'd51: q = 32'hc3c35e9d;
	8'd52: q = 32'h18182830;
	8'd53: q = 32'h9696a137;
	8'd54: q = 32'h5050f0a;
	8'd55: q = 32'h9a9ab52f;
	8'd56: q = 32'h707090e;
	8'd57: q = 32'h12123624;
	8'd58: q = 32'h80809b1b;
	8'd59: q = 32'he2e23ddf;
	8'd60: q = 32'hebeb26cd;
	8'd61: q = 32'h2727694e;
	8'd62: q = 32'hb2b2cd7f;
	8'd63: q = 32'h75759fea;
	8'd64: q = 32'h9091b12;
	8'd65: q = 32'h83839e1d;
	8'd66: q = 32'h2c2c7458;
	8'd67: q = 32'h1a1a2e34;
	8'd68: q = 32'h1b1b2d36;
	8'd69: q = 32'h6e6eb2dc;
	8'd70: q = 32'h5a5aeeb4;
	8'd71: q = 32'ha0a0fb5b;
	8'd72: q = 32'h5252f6a4;
	8'd73: q = 32'h3b3b4d76;
	8'd74: q = 32'hd6d661b7;
	8'd75: q = 32'hb3b3ce7d;
	8'd76: q = 32'h29297b52;
	8'd77: q = 32'he3e33edd;
	8'd78: q = 32'h2f2f715e;
	8'd79: q = 32'h84849713;
	8'd80: q = 32'h5353f5a6;
	8'd81: q = 32'hd1d168b9;
	8'd82: q = 32'h0;
	8'd83: q = 32'heded2cc1;
	8'd84: q = 32'h20206040;
	8'd85: q = 32'hfcfc1fe3;
	8'd86: q = 32'hb1b1c879;
	8'd87: q = 32'h5b5bedb6;
	8'd88: q = 32'h6a6abed4;
	8'd89: q = 32'hcbcb468d;
	8'd90: q = 32'hbebed967;
	8'd91: q = 32'h39394b72;
	8'd92: q = 32'h4a4ade94;
	8'd93: q = 32'h4c4cd498;
	8'd94: q = 32'h5858e8b0;
	8'd95: q = 32'hcfcf4a85;
	8'd96: q = 32'hd0d06bbb;
	8'd97: q = 32'hefef2ac5;
	8'd98: q = 32'haaaae54f;
	8'd99: q = 32'hfbfb16ed;
	8'd100: q = 32'h4343c586;
	8'd101: q = 32'h4d4dd79a;
	8'd102: q = 32'h33335566;
	8'd103: q = 32'h85859411;
	8'd104: q = 32'h4545cf8a;
	8'd105: q = 32'hf9f910e9;
	8'd106: q = 32'h2020604;
	8'd107: q = 32'h7f7f81fe;
	8'd108: q = 32'h5050f0a0;
	8'd109: q = 32'h3c3c4478;
	8'd110: q = 32'h9f9fba25;
	8'd111: q = 32'ha8a8e34b;
	8'd112: q = 32'h5151f3a2;
	8'd113: q = 32'ha3a3fe5d;
	8'd114: q = 32'h4040c080;
	8'd115: q = 32'h8f8f8a05;
	8'd116: q = 32'h9292ad3f;
	8'd117: q = 32'h9d9dbc21;
	8'd118: q = 32'h38384870;
	8'd119: q = 32'hf5f504f1;
	8'd120: q = 32'hbcbcdf63;
	8'd121: q = 32'hb6b6c177;
	8'd122: q = 32'hdada75af;
	8'd123: q = 32'h21216342;
	8'd124: q = 32'h10103020;
	8'd125: q = 32'hffff1ae5;
	8'd126: q = 32'hf3f30efd;
	8'd127: q = 32'hd2d26dbf;
	8'd128: q = 32'hcdcd4c81;
	8'd129: q = 32'hc0c1418;
	8'd130: q = 32'h13133526;
	8'd131: q = 32'hecec2fc3;
	8'd132: q = 32'h5f5fe1be;
	8'd133: q = 32'h9797a235;
	8'd134: q = 32'h4444cc88;
	8'd135: q = 32'h1717392e;
	8'd136: q = 32'hc4c45793;
	8'd137: q = 32'ha7a7f255;
	8'd138: q = 32'h7e7e82fc;
	8'd139: q = 32'h3d3d477a;
	8'd140: q = 32'h6464acc8;
	8'd141: q = 32'h5d5de7ba;
	8'd142: q = 32'h19192b32;
	8'd143: q = 32'h737395e6;
	8'd144: q = 32'h6060a0c0;
	8'd145: q = 32'h81819819;
	8'd146: q = 32'h4f4fd19e;
	8'd147: q = 32'hdcdc7fa3;
	8'd148: q = 32'h22226644;
	8'd149: q = 32'h2a2a7e54;
	8'd150: q = 32'h9090ab3b;
	8'd151: q = 32'h8888830b;
	8'd152: q = 32'h4646ca8c;
	8'd153: q = 32'heeee29c7;
	8'd154: q = 32'hb8b8d36b;
	8'd155: q = 32'h14143c28;
	8'd156: q = 32'hdede79a7;
	8'd157: q = 32'h5e5ee2bc;
	8'd158: q = 32'hb0b1d16;
	8'd159: q = 32'hdbdb76ad;
	8'd160: q = 32'he0e03bdb;
	8'd161: q = 32'h32325664;
	8'd162: q = 32'h3a3a4e74;
	8'd163: q = 32'ha0a1e14;
	8'd164: q = 32'h4949db92;
	8'd165: q = 32'h6060a0c;
	8'd166: q = 32'h24246c48;
	8'd167: q = 32'h5c5ce4b8;
	8'd168: q = 32'hc2c25d9f;
	8'd169: q = 32'hd3d36ebd;
	8'd170: q = 32'hacacef43;
	8'd171: q = 32'h6262a6c4;
	8'd172: q = 32'h9191a839;
	8'd173: q = 32'h9595a431;
	8'd174: q = 32'he4e437d3;
	8'd175: q = 32'h79798bf2;
	8'd176: q = 32'he7e732d5;
	8'd177: q = 32'hc8c8438b;
	8'd178: q = 32'h3737596e;
	8'd179: q = 32'h6d6db7da;
	8'd180: q = 32'h8d8d8c01;
	8'd181: q = 32'hd5d564b1;
	8'd182: q = 32'h4e4ed29c;
	8'd183: q = 32'ha9a9e049;
	8'd184: q = 32'h6c6cb4d8;
	8'd185: q = 32'h5656faac;
	8'd186: q = 32'hf4f407f3;
	8'd187: q = 32'heaea25cf;
	8'd188: q = 32'h6565afca;
	8'd189: q = 32'h7a7a8ef4;
	8'd190: q = 32'haeaee947;
	8'd191: q = 32'h8081810;
	8'd192: q = 32'hbabad56f;
	8'd193: q = 32'h787888f0;
	8'd194: q = 32'h25256f4a;
	8'd195: q = 32'h2e2e725c;
	8'd196: q = 32'h1c1c2438;
	8'd197: q = 32'ha6a6f157;
	8'd198: q = 32'hb4b4c773;
	8'd199: q = 32'hc6c65197;
	8'd200: q = 32'he8e823cb;
	8'd201: q = 32'hdddd7ca1;
	8'd202: q = 32'h74749ce8;
	8'd203: q = 32'h1f1f213e;
	8'd204: q = 32'h4b4bdd96;
	8'd205: q = 32'hbdbddc61;
	8'd206: q = 32'h8b8b860d;
	8'd207: q = 32'h8a8a850f;
	8'd208: q = 32'h707090e0;
	8'd209: q = 32'h3e3e427c;
	8'd210: q = 32'hb5b5c471;
	8'd211: q = 32'h6666aacc;
	8'd212: q = 32'h4848d890;
	8'd213: q = 32'h3030506;
	8'd214: q = 32'hf6f601f7;
	8'd215: q = 32'he0e121c;
	8'd216: q = 32'h6161a3c2;
	8'd217: q = 32'h35355f6a;
	8'd218: q = 32'h5757f9ae;
	8'd219: q = 32'hb9b9d069;
	8'd220: q = 32'h86869117;
	8'd221: q = 32'hc1c15899;
	8'd222: q = 32'h1d1d273a;
	8'd223: q = 32'h9e9eb927;
	8'd224: q = 32'he1e138d9;
	8'd225: q = 32'hf8f813eb;
	8'd226: q = 32'h9898b32b;
	8'd227: q = 32'h11113322;
	8'd228: q = 32'h6969bbd2;
	8'd229: q = 32'hd9d970a9;
	8'd230: q = 32'h8e8e8907;
	8'd231: q = 32'h9494a733;
	8'd232: q = 32'h9b9bb62d;
	8'd233: q = 32'h1e1e223c;
	8'd234: q = 32'h87879215;
	8'd235: q = 32'he9e920c9;
	8'd236: q = 32'hcece4987;
	8'd237: q = 32'h5555ffaa;
	8'd238: q = 32'h28287850;
	8'd239: q = 32'hdfdf7aa5;
	8'd240: q = 32'h8c8c8f03;
	8'd241: q = 32'ha1a1f859;
	8'd242: q = 32'h89898009;
	8'd243: q = 32'hd0d171a;
	8'd244: q = 32'hbfbfda65;
	8'd245: q = 32'he6e631d7;
	8'd246: q = 32'h4242c684;
	8'd247: q = 32'h6868b8d0;
	8'd248: q = 32'h4141c382;
	8'd249: q = 32'h9999b029;
	8'd250: q = 32'h2d2d775a;
	8'd251: q = 32'hf0f111e;
	8'd252: q = 32'hb0b0cb7b;
	8'd253: q = 32'h5454fca8;
	8'd254: q = 32'hbbbbd66d;
	8'd255: q = 32'h16163a2c;

     endcase // case (a)
endmodule

