module tboxe1(input wire clk,
              input wire [7:0] a,
              output reg [31:0] q);

   always @(posedge clk)
     case (a)
	8'd0: q = 32'ha5c66363;
	8'd1: q = 32'h84f87c7c;
	8'd2: q = 32'h99ee7777;
	8'd3: q = 32'h8df67b7b;
	8'd4: q = 32'hdfff2f2;
	8'd5: q = 32'hbdd66b6b;
	8'd6: q = 32'hb1de6f6f;
	8'd7: q = 32'h5491c5c5;
	8'd8: q = 32'h50603030;
	8'd9: q = 32'h3020101;
	8'd10: q = 32'ha9ce6767;
	8'd11: q = 32'h7d562b2b;
	8'd12: q = 32'h19e7fefe;
	8'd13: q = 32'h62b5d7d7;
	8'd14: q = 32'he64dabab;
	8'd15: q = 32'h9aec7676;
	8'd16: q = 32'h458fcaca;
	8'd17: q = 32'h9d1f8282;
	8'd18: q = 32'h4089c9c9;
	8'd19: q = 32'h87fa7d7d;
	8'd20: q = 32'h15effafa;
	8'd21: q = 32'hebb25959;
	8'd22: q = 32'hc98e4747;
	8'd23: q = 32'hbfbf0f0;
	8'd24: q = 32'hec41adad;
	8'd25: q = 32'h67b3d4d4;
	8'd26: q = 32'hfd5fa2a2;
	8'd27: q = 32'hea45afaf;
	8'd28: q = 32'hbf239c9c;
	8'd29: q = 32'hf753a4a4;
	8'd30: q = 32'h96e47272;
	8'd31: q = 32'h5b9bc0c0;
	8'd32: q = 32'hc275b7b7;
	8'd33: q = 32'h1ce1fdfd;
	8'd34: q = 32'hae3d9393;
	8'd35: q = 32'h6a4c2626;
	8'd36: q = 32'h5a6c3636;
	8'd37: q = 32'h417e3f3f;
	8'd38: q = 32'h2f5f7f7;
	8'd39: q = 32'h4f83cccc;
	8'd40: q = 32'h5c683434;
	8'd41: q = 32'hf451a5a5;
	8'd42: q = 32'h34d1e5e5;
	8'd43: q = 32'h8f9f1f1;
	8'd44: q = 32'h93e27171;
	8'd45: q = 32'h73abd8d8;
	8'd46: q = 32'h53623131;
	8'd47: q = 32'h3f2a1515;
	8'd48: q = 32'hc080404;
	8'd49: q = 32'h5295c7c7;
	8'd50: q = 32'h65462323;
	8'd51: q = 32'h5e9dc3c3;
	8'd52: q = 32'h28301818;
	8'd53: q = 32'ha1379696;
	8'd54: q = 32'hf0a0505;
	8'd55: q = 32'hb52f9a9a;
	8'd56: q = 32'h90e0707;
	8'd57: q = 32'h36241212;
	8'd58: q = 32'h9b1b8080;
	8'd59: q = 32'h3ddfe2e2;
	8'd60: q = 32'h26cdebeb;
	8'd61: q = 32'h694e2727;
	8'd62: q = 32'hcd7fb2b2;
	8'd63: q = 32'h9fea7575;
	8'd64: q = 32'h1b120909;
	8'd65: q = 32'h9e1d8383;
	8'd66: q = 32'h74582c2c;
	8'd67: q = 32'h2e341a1a;
	8'd68: q = 32'h2d361b1b;
	8'd69: q = 32'hb2dc6e6e;
	8'd70: q = 32'heeb45a5a;
	8'd71: q = 32'hfb5ba0a0;
	8'd72: q = 32'hf6a45252;
	8'd73: q = 32'h4d763b3b;
	8'd74: q = 32'h61b7d6d6;
	8'd75: q = 32'hce7db3b3;
	8'd76: q = 32'h7b522929;
	8'd77: q = 32'h3edde3e3;
	8'd78: q = 32'h715e2f2f;
	8'd79: q = 32'h97138484;
	8'd80: q = 32'hf5a65353;
	8'd81: q = 32'h68b9d1d1;
	8'd82: q = 32'h0;
	8'd83: q = 32'h2cc1eded;
	8'd84: q = 32'h60402020;
	8'd85: q = 32'h1fe3fcfc;
	8'd86: q = 32'hc879b1b1;
	8'd87: q = 32'hedb65b5b;
	8'd88: q = 32'hbed46a6a;
	8'd89: q = 32'h468dcbcb;
	8'd90: q = 32'hd967bebe;
	8'd91: q = 32'h4b723939;
	8'd92: q = 32'hde944a4a;
	8'd93: q = 32'hd4984c4c;
	8'd94: q = 32'he8b05858;
	8'd95: q = 32'h4a85cfcf;
	8'd96: q = 32'h6bbbd0d0;
	8'd97: q = 32'h2ac5efef;
	8'd98: q = 32'he54faaaa;
	8'd99: q = 32'h16edfbfb;
	8'd100: q = 32'hc5864343;
	8'd101: q = 32'hd79a4d4d;
	8'd102: q = 32'h55663333;
	8'd103: q = 32'h94118585;
	8'd104: q = 32'hcf8a4545;
	8'd105: q = 32'h10e9f9f9;
	8'd106: q = 32'h6040202;
	8'd107: q = 32'h81fe7f7f;
	8'd108: q = 32'hf0a05050;
	8'd109: q = 32'h44783c3c;
	8'd110: q = 32'hba259f9f;
	8'd111: q = 32'he34ba8a8;
	8'd112: q = 32'hf3a25151;
	8'd113: q = 32'hfe5da3a3;
	8'd114: q = 32'hc0804040;
	8'd115: q = 32'h8a058f8f;
	8'd116: q = 32'had3f9292;
	8'd117: q = 32'hbc219d9d;
	8'd118: q = 32'h48703838;
	8'd119: q = 32'h4f1f5f5;
	8'd120: q = 32'hdf63bcbc;
	8'd121: q = 32'hc177b6b6;
	8'd122: q = 32'h75afdada;
	8'd123: q = 32'h63422121;
	8'd124: q = 32'h30201010;
	8'd125: q = 32'h1ae5ffff;
	8'd126: q = 32'hefdf3f3;
	8'd127: q = 32'h6dbfd2d2;
	8'd128: q = 32'h4c81cdcd;
	8'd129: q = 32'h14180c0c;
	8'd130: q = 32'h35261313;
	8'd131: q = 32'h2fc3ecec;
	8'd132: q = 32'he1be5f5f;
	8'd133: q = 32'ha2359797;
	8'd134: q = 32'hcc884444;
	8'd135: q = 32'h392e1717;
	8'd136: q = 32'h5793c4c4;
	8'd137: q = 32'hf255a7a7;
	8'd138: q = 32'h82fc7e7e;
	8'd139: q = 32'h477a3d3d;
	8'd140: q = 32'hacc86464;
	8'd141: q = 32'he7ba5d5d;
	8'd142: q = 32'h2b321919;
	8'd143: q = 32'h95e67373;
	8'd144: q = 32'ha0c06060;
	8'd145: q = 32'h98198181;
	8'd146: q = 32'hd19e4f4f;
	8'd147: q = 32'h7fa3dcdc;
	8'd148: q = 32'h66442222;
	8'd149: q = 32'h7e542a2a;
	8'd150: q = 32'hab3b9090;
	8'd151: q = 32'h830b8888;
	8'd152: q = 32'hca8c4646;
	8'd153: q = 32'h29c7eeee;
	8'd154: q = 32'hd36bb8b8;
	8'd155: q = 32'h3c281414;
	8'd156: q = 32'h79a7dede;
	8'd157: q = 32'he2bc5e5e;
	8'd158: q = 32'h1d160b0b;
	8'd159: q = 32'h76addbdb;
	8'd160: q = 32'h3bdbe0e0;
	8'd161: q = 32'h56643232;
	8'd162: q = 32'h4e743a3a;
	8'd163: q = 32'h1e140a0a;
	8'd164: q = 32'hdb924949;
	8'd165: q = 32'ha0c0606;
	8'd166: q = 32'h6c482424;
	8'd167: q = 32'he4b85c5c;
	8'd168: q = 32'h5d9fc2c2;
	8'd169: q = 32'h6ebdd3d3;
	8'd170: q = 32'hef43acac;
	8'd171: q = 32'ha6c46262;
	8'd172: q = 32'ha8399191;
	8'd173: q = 32'ha4319595;
	8'd174: q = 32'h37d3e4e4;
	8'd175: q = 32'h8bf27979;
	8'd176: q = 32'h32d5e7e7;
	8'd177: q = 32'h438bc8c8;
	8'd178: q = 32'h596e3737;
	8'd179: q = 32'hb7da6d6d;
	8'd180: q = 32'h8c018d8d;
	8'd181: q = 32'h64b1d5d5;
	8'd182: q = 32'hd29c4e4e;
	8'd183: q = 32'he049a9a9;
	8'd184: q = 32'hb4d86c6c;
	8'd185: q = 32'hfaac5656;
	8'd186: q = 32'h7f3f4f4;
	8'd187: q = 32'h25cfeaea;
	8'd188: q = 32'hafca6565;
	8'd189: q = 32'h8ef47a7a;
	8'd190: q = 32'he947aeae;
	8'd191: q = 32'h18100808;
	8'd192: q = 32'hd56fbaba;
	8'd193: q = 32'h88f07878;
	8'd194: q = 32'h6f4a2525;
	8'd195: q = 32'h725c2e2e;
	8'd196: q = 32'h24381c1c;
	8'd197: q = 32'hf157a6a6;
	8'd198: q = 32'hc773b4b4;
	8'd199: q = 32'h5197c6c6;
	8'd200: q = 32'h23cbe8e8;
	8'd201: q = 32'h7ca1dddd;
	8'd202: q = 32'h9ce87474;
	8'd203: q = 32'h213e1f1f;
	8'd204: q = 32'hdd964b4b;
	8'd205: q = 32'hdc61bdbd;
	8'd206: q = 32'h860d8b8b;
	8'd207: q = 32'h850f8a8a;
	8'd208: q = 32'h90e07070;
	8'd209: q = 32'h427c3e3e;
	8'd210: q = 32'hc471b5b5;
	8'd211: q = 32'haacc6666;
	8'd212: q = 32'hd8904848;
	8'd213: q = 32'h5060303;
	8'd214: q = 32'h1f7f6f6;
	8'd215: q = 32'h121c0e0e;
	8'd216: q = 32'ha3c26161;
	8'd217: q = 32'h5f6a3535;
	8'd218: q = 32'hf9ae5757;
	8'd219: q = 32'hd069b9b9;
	8'd220: q = 32'h91178686;
	8'd221: q = 32'h5899c1c1;
	8'd222: q = 32'h273a1d1d;
	8'd223: q = 32'hb9279e9e;
	8'd224: q = 32'h38d9e1e1;
	8'd225: q = 32'h13ebf8f8;
	8'd226: q = 32'hb32b9898;
	8'd227: q = 32'h33221111;
	8'd228: q = 32'hbbd26969;
	8'd229: q = 32'h70a9d9d9;
	8'd230: q = 32'h89078e8e;
	8'd231: q = 32'ha7339494;
	8'd232: q = 32'hb62d9b9b;
	8'd233: q = 32'h223c1e1e;
	8'd234: q = 32'h92158787;
	8'd235: q = 32'h20c9e9e9;
	8'd236: q = 32'h4987cece;
	8'd237: q = 32'hffaa5555;
	8'd238: q = 32'h78502828;
	8'd239: q = 32'h7aa5dfdf;
	8'd240: q = 32'h8f038c8c;
	8'd241: q = 32'hf859a1a1;
	8'd242: q = 32'h80098989;
	8'd243: q = 32'h171a0d0d;
	8'd244: q = 32'hda65bfbf;
	8'd245: q = 32'h31d7e6e6;
	8'd246: q = 32'hc6844242;
	8'd247: q = 32'hb8d06868;
	8'd248: q = 32'hc3824141;
	8'd249: q = 32'hb0299999;
	8'd250: q = 32'h775a2d2d;
	8'd251: q = 32'h111e0f0f;
	8'd252: q = 32'hcb7bb0b0;
	8'd253: q = 32'hfca85454;
	8'd254: q = 32'hd66dbbbb;
	8'd255: q = 32'h3a2c1616;

     endcase // case (a)
endmodule

