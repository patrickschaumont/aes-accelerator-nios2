module tboxe0(input wire clk,
              input wire [7:0] a,
              output reg [31:0] q);

   always @(posedge clk)
     case (a)
	8'd0: q = 32'hc66363a5;
	8'd1: q = 32'hf87c7c84;
	8'd2: q = 32'hee777799;
	8'd3: q = 32'hf67b7b8d;
	8'd4: q = 32'hfff2f20d;
	8'd5: q = 32'hd66b6bbd;
	8'd6: q = 32'hde6f6fb1;
	8'd7: q = 32'h91c5c554;
	8'd8: q = 32'h60303050;
	8'd9: q = 32'h2010103;
	8'd10: q = 32'hce6767a9;
	8'd11: q = 32'h562b2b7d;
	8'd12: q = 32'he7fefe19;
	8'd13: q = 32'hb5d7d762;
	8'd14: q = 32'h4dababe6;
	8'd15: q = 32'hec76769a;
	8'd16: q = 32'h8fcaca45;
	8'd17: q = 32'h1f82829d;
	8'd18: q = 32'h89c9c940;
	8'd19: q = 32'hfa7d7d87;
	8'd20: q = 32'heffafa15;
	8'd21: q = 32'hb25959eb;
	8'd22: q = 32'h8e4747c9;
	8'd23: q = 32'hfbf0f00b;
	8'd24: q = 32'h41adadec;
	8'd25: q = 32'hb3d4d467;
	8'd26: q = 32'h5fa2a2fd;
	8'd27: q = 32'h45afafea;
	8'd28: q = 32'h239c9cbf;
	8'd29: q = 32'h53a4a4f7;
	8'd30: q = 32'he4727296;
	8'd31: q = 32'h9bc0c05b;
	8'd32: q = 32'h75b7b7c2;
	8'd33: q = 32'he1fdfd1c;
	8'd34: q = 32'h3d9393ae;
	8'd35: q = 32'h4c26266a;
	8'd36: q = 32'h6c36365a;
	8'd37: q = 32'h7e3f3f41;
	8'd38: q = 32'hf5f7f702;
	8'd39: q = 32'h83cccc4f;
	8'd40: q = 32'h6834345c;
	8'd41: q = 32'h51a5a5f4;
	8'd42: q = 32'hd1e5e534;
	8'd43: q = 32'hf9f1f108;
	8'd44: q = 32'he2717193;
	8'd45: q = 32'habd8d873;
	8'd46: q = 32'h62313153;
	8'd47: q = 32'h2a15153f;
	8'd48: q = 32'h804040c;
	8'd49: q = 32'h95c7c752;
	8'd50: q = 32'h46232365;
	8'd51: q = 32'h9dc3c35e;
	8'd52: q = 32'h30181828;
	8'd53: q = 32'h379696a1;
	8'd54: q = 32'ha05050f;
	8'd55: q = 32'h2f9a9ab5;
	8'd56: q = 32'he070709;
	8'd57: q = 32'h24121236;
	8'd58: q = 32'h1b80809b;
	8'd59: q = 32'hdfe2e23d;
	8'd60: q = 32'hcdebeb26;
	8'd61: q = 32'h4e272769;
	8'd62: q = 32'h7fb2b2cd;
	8'd63: q = 32'hea75759f;
	8'd64: q = 32'h1209091b;
	8'd65: q = 32'h1d83839e;
	8'd66: q = 32'h582c2c74;
	8'd67: q = 32'h341a1a2e;
	8'd68: q = 32'h361b1b2d;
	8'd69: q = 32'hdc6e6eb2;
	8'd70: q = 32'hb45a5aee;
	8'd71: q = 32'h5ba0a0fb;
	8'd72: q = 32'ha45252f6;
	8'd73: q = 32'h763b3b4d;
	8'd74: q = 32'hb7d6d661;
	8'd75: q = 32'h7db3b3ce;
	8'd76: q = 32'h5229297b;
	8'd77: q = 32'hdde3e33e;
	8'd78: q = 32'h5e2f2f71;
	8'd79: q = 32'h13848497;
	8'd80: q = 32'ha65353f5;
	8'd81: q = 32'hb9d1d168;
	8'd82: q = 32'h0;
	8'd83: q = 32'hc1eded2c;
	8'd84: q = 32'h40202060;
	8'd85: q = 32'he3fcfc1f;
	8'd86: q = 32'h79b1b1c8;
	8'd87: q = 32'hb65b5bed;
	8'd88: q = 32'hd46a6abe;
	8'd89: q = 32'h8dcbcb46;
	8'd90: q = 32'h67bebed9;
	8'd91: q = 32'h7239394b;
	8'd92: q = 32'h944a4ade;
	8'd93: q = 32'h984c4cd4;
	8'd94: q = 32'hb05858e8;
	8'd95: q = 32'h85cfcf4a;
	8'd96: q = 32'hbbd0d06b;
	8'd97: q = 32'hc5efef2a;
	8'd98: q = 32'h4faaaae5;
	8'd99: q = 32'hedfbfb16;
	8'd100: q = 32'h864343c5;
	8'd101: q = 32'h9a4d4dd7;
	8'd102: q = 32'h66333355;
	8'd103: q = 32'h11858594;
	8'd104: q = 32'h8a4545cf;
	8'd105: q = 32'he9f9f910;
	8'd106: q = 32'h4020206;
	8'd107: q = 32'hfe7f7f81;
	8'd108: q = 32'ha05050f0;
	8'd109: q = 32'h783c3c44;
	8'd110: q = 32'h259f9fba;
	8'd111: q = 32'h4ba8a8e3;
	8'd112: q = 32'ha25151f3;
	8'd113: q = 32'h5da3a3fe;
	8'd114: q = 32'h804040c0;
	8'd115: q = 32'h58f8f8a;
	8'd116: q = 32'h3f9292ad;
	8'd117: q = 32'h219d9dbc;
	8'd118: q = 32'h70383848;
	8'd119: q = 32'hf1f5f504;
	8'd120: q = 32'h63bcbcdf;
	8'd121: q = 32'h77b6b6c1;
	8'd122: q = 32'hafdada75;
	8'd123: q = 32'h42212163;
	8'd124: q = 32'h20101030;
	8'd125: q = 32'he5ffff1a;
	8'd126: q = 32'hfdf3f30e;
	8'd127: q = 32'hbfd2d26d;
	8'd128: q = 32'h81cdcd4c;
	8'd129: q = 32'h180c0c14;
	8'd130: q = 32'h26131335;
	8'd131: q = 32'hc3ecec2f;
	8'd132: q = 32'hbe5f5fe1;
	8'd133: q = 32'h359797a2;
	8'd134: q = 32'h884444cc;
	8'd135: q = 32'h2e171739;
	8'd136: q = 32'h93c4c457;
	8'd137: q = 32'h55a7a7f2;
	8'd138: q = 32'hfc7e7e82;
	8'd139: q = 32'h7a3d3d47;
	8'd140: q = 32'hc86464ac;
	8'd141: q = 32'hba5d5de7;
	8'd142: q = 32'h3219192b;
	8'd143: q = 32'he6737395;
	8'd144: q = 32'hc06060a0;
	8'd145: q = 32'h19818198;
	8'd146: q = 32'h9e4f4fd1;
	8'd147: q = 32'ha3dcdc7f;
	8'd148: q = 32'h44222266;
	8'd149: q = 32'h542a2a7e;
	8'd150: q = 32'h3b9090ab;
	8'd151: q = 32'hb888883;
	8'd152: q = 32'h8c4646ca;
	8'd153: q = 32'hc7eeee29;
	8'd154: q = 32'h6bb8b8d3;
	8'd155: q = 32'h2814143c;
	8'd156: q = 32'ha7dede79;
	8'd157: q = 32'hbc5e5ee2;
	8'd158: q = 32'h160b0b1d;
	8'd159: q = 32'haddbdb76;
	8'd160: q = 32'hdbe0e03b;
	8'd161: q = 32'h64323256;
	8'd162: q = 32'h743a3a4e;
	8'd163: q = 32'h140a0a1e;
	8'd164: q = 32'h924949db;
	8'd165: q = 32'hc06060a;
	8'd166: q = 32'h4824246c;
	8'd167: q = 32'hb85c5ce4;
	8'd168: q = 32'h9fc2c25d;
	8'd169: q = 32'hbdd3d36e;
	8'd170: q = 32'h43acacef;
	8'd171: q = 32'hc46262a6;
	8'd172: q = 32'h399191a8;
	8'd173: q = 32'h319595a4;
	8'd174: q = 32'hd3e4e437;
	8'd175: q = 32'hf279798b;
	8'd176: q = 32'hd5e7e732;
	8'd177: q = 32'h8bc8c843;
	8'd178: q = 32'h6e373759;
	8'd179: q = 32'hda6d6db7;
	8'd180: q = 32'h18d8d8c;
	8'd181: q = 32'hb1d5d564;
	8'd182: q = 32'h9c4e4ed2;
	8'd183: q = 32'h49a9a9e0;
	8'd184: q = 32'hd86c6cb4;
	8'd185: q = 32'hac5656fa;
	8'd186: q = 32'hf3f4f407;
	8'd187: q = 32'hcfeaea25;
	8'd188: q = 32'hca6565af;
	8'd189: q = 32'hf47a7a8e;
	8'd190: q = 32'h47aeaee9;
	8'd191: q = 32'h10080818;
	8'd192: q = 32'h6fbabad5;
	8'd193: q = 32'hf0787888;
	8'd194: q = 32'h4a25256f;
	8'd195: q = 32'h5c2e2e72;
	8'd196: q = 32'h381c1c24;
	8'd197: q = 32'h57a6a6f1;
	8'd198: q = 32'h73b4b4c7;
	8'd199: q = 32'h97c6c651;
	8'd200: q = 32'hcbe8e823;
	8'd201: q = 32'ha1dddd7c;
	8'd202: q = 32'he874749c;
	8'd203: q = 32'h3e1f1f21;
	8'd204: q = 32'h964b4bdd;
	8'd205: q = 32'h61bdbddc;
	8'd206: q = 32'hd8b8b86;
	8'd207: q = 32'hf8a8a85;
	8'd208: q = 32'he0707090;
	8'd209: q = 32'h7c3e3e42;
	8'd210: q = 32'h71b5b5c4;
	8'd211: q = 32'hcc6666aa;
	8'd212: q = 32'h904848d8;
	8'd213: q = 32'h6030305;
	8'd214: q = 32'hf7f6f601;
	8'd215: q = 32'h1c0e0e12;
	8'd216: q = 32'hc26161a3;
	8'd217: q = 32'h6a35355f;
	8'd218: q = 32'hae5757f9;
	8'd219: q = 32'h69b9b9d0;
	8'd220: q = 32'h17868691;
	8'd221: q = 32'h99c1c158;
	8'd222: q = 32'h3a1d1d27;
	8'd223: q = 32'h279e9eb9;
	8'd224: q = 32'hd9e1e138;
	8'd225: q = 32'hebf8f813;
	8'd226: q = 32'h2b9898b3;
	8'd227: q = 32'h22111133;
	8'd228: q = 32'hd26969bb;
	8'd229: q = 32'ha9d9d970;
	8'd230: q = 32'h78e8e89;
	8'd231: q = 32'h339494a7;
	8'd232: q = 32'h2d9b9bb6;
	8'd233: q = 32'h3c1e1e22;
	8'd234: q = 32'h15878792;
	8'd235: q = 32'hc9e9e920;
	8'd236: q = 32'h87cece49;
	8'd237: q = 32'haa5555ff;
	8'd238: q = 32'h50282878;
	8'd239: q = 32'ha5dfdf7a;
	8'd240: q = 32'h38c8c8f;
	8'd241: q = 32'h59a1a1f8;
	8'd242: q = 32'h9898980;
	8'd243: q = 32'h1a0d0d17;
	8'd244: q = 32'h65bfbfda;
	8'd245: q = 32'hd7e6e631;
	8'd246: q = 32'h844242c6;
	8'd247: q = 32'hd06868b8;
	8'd248: q = 32'h824141c3;
	8'd249: q = 32'h299999b0;
	8'd250: q = 32'h5a2d2d77;
	8'd251: q = 32'h1e0f0f11;
	8'd252: q = 32'h7bb0b0cb;
	8'd253: q = 32'ha85454fc;
	8'd254: q = 32'h6dbbbbd6;
	8'd255: q = 32'h2c16163a;

     endcase // case (a)
endmodule

