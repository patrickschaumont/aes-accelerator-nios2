module tboxd3(input wire clk,
              input wire [7:0] a,
              output reg [31:0] q);

   always @(posedge clk)
     case (a)
	8'd0: q = 32'hf4a75051;
	8'd1: q = 32'h4165537e;
	8'd2: q = 32'h17a4c31a;
	8'd3: q = 32'h275e963a;
	8'd4: q = 32'hab6bcb3b;
	8'd5: q = 32'h9d45f11f;
	8'd6: q = 32'hfa58abac;
	8'd7: q = 32'he303934b;
	8'd8: q = 32'h30fa5520;
	8'd9: q = 32'h766df6ad;
	8'd10: q = 32'hcc769188;
	8'd11: q = 32'h24c25f5;
	8'd12: q = 32'he5d7fc4f;
	8'd13: q = 32'h2acbd7c5;
	8'd14: q = 32'h35448026;
	8'd15: q = 32'h62a38fb5;
	8'd16: q = 32'hb15a49de;
	8'd17: q = 32'hba1b6725;
	8'd18: q = 32'hea0e9845;
	8'd19: q = 32'hfec0e15d;
	8'd20: q = 32'h2f7502c3;
	8'd21: q = 32'h4cf01281;
	8'd22: q = 32'h4697a38d;
	8'd23: q = 32'hd3f9c66b;
	8'd24: q = 32'h8f5fe703;
	8'd25: q = 32'h929c9515;
	8'd26: q = 32'h6d7aebbf;
	8'd27: q = 32'h5259da95;
	8'd28: q = 32'hbe832dd4;
	8'd29: q = 32'h7421d358;
	8'd30: q = 32'he0692949;
	8'd31: q = 32'hc9c8448e;
	8'd32: q = 32'hc2896a75;
	8'd33: q = 32'h8e7978f4;
	8'd34: q = 32'h583e6b99;
	8'd35: q = 32'hb971dd27;
	8'd36: q = 32'he14fb6be;
	8'd37: q = 32'h88ad17f0;
	8'd38: q = 32'h20ac66c9;
	8'd39: q = 32'hce3ab47d;
	8'd40: q = 32'hdf4a1863;
	8'd41: q = 32'h1a3182e5;
	8'd42: q = 32'h51336097;
	8'd43: q = 32'h537f4562;
	8'd44: q = 32'h6477e0b1;
	8'd45: q = 32'h6bae84bb;
	8'd46: q = 32'h81a01cfe;
	8'd47: q = 32'h82b94f9;
	8'd48: q = 32'h48685870;
	8'd49: q = 32'h45fd198f;
	8'd50: q = 32'hde6c8794;
	8'd51: q = 32'h7bf8b752;
	8'd52: q = 32'h73d323ab;
	8'd53: q = 32'h4b02e272;
	8'd54: q = 32'h1f8f57e3;
	8'd55: q = 32'h55ab2a66;
	8'd56: q = 32'heb2807b2;
	8'd57: q = 32'hb5c2032f;
	8'd58: q = 32'hc57b9a86;
	8'd59: q = 32'h3708a5d3;
	8'd60: q = 32'h2887f230;
	8'd61: q = 32'hbfa5b223;
	8'd62: q = 32'h36aba02;
	8'd63: q = 32'h16825ced;
	8'd64: q = 32'hcf1c2b8a;
	8'd65: q = 32'h79b492a7;
	8'd66: q = 32'h7f2f0f3;
	8'd67: q = 32'h69e2a14e;
	8'd68: q = 32'hdaf4cd65;
	8'd69: q = 32'h5bed506;
	8'd70: q = 32'h34621fd1;
	8'd71: q = 32'ha6fe8ac4;
	8'd72: q = 32'h2e539d34;
	8'd73: q = 32'hf355a0a2;
	8'd74: q = 32'h8ae13205;
	8'd75: q = 32'hf6eb75a4;
	8'd76: q = 32'h83ec390b;
	8'd77: q = 32'h60efaa40;
	8'd78: q = 32'h719f065e;
	8'd79: q = 32'h6e1051bd;
	8'd80: q = 32'h218af93e;
	8'd81: q = 32'hdd063d96;
	8'd82: q = 32'h3e05aedd;
	8'd83: q = 32'he6bd464d;
	8'd84: q = 32'h548db591;
	8'd85: q = 32'hc45d0571;
	8'd86: q = 32'h6d46f04;
	8'd87: q = 32'h5015ff60;
	8'd88: q = 32'h98fb2419;
	8'd89: q = 32'hbde997d6;
	8'd90: q = 32'h4043cc89;
	8'd91: q = 32'hd99e7767;
	8'd92: q = 32'he842bdb0;
	8'd93: q = 32'h898b8807;
	8'd94: q = 32'h195b38e7;
	8'd95: q = 32'hc8eedb79;
	8'd96: q = 32'h7c0a47a1;
	8'd97: q = 32'h420fe97c;
	8'd98: q = 32'h841ec9f8;
	8'd99: q = 32'h0;
	8'd100: q = 32'h80868309;
	8'd101: q = 32'h2bed4832;
	8'd102: q = 32'h1170ac1e;
	8'd103: q = 32'h5a724e6c;
	8'd104: q = 32'hefffbfd;
	8'd105: q = 32'h8538560f;
	8'd106: q = 32'haed51e3d;
	8'd107: q = 32'h2d392736;
	8'd108: q = 32'hfd9640a;
	8'd109: q = 32'h5ca62168;
	8'd110: q = 32'h5b54d19b;
	8'd111: q = 32'h362e3a24;
	8'd112: q = 32'ha67b10c;
	8'd113: q = 32'h57e70f93;
	8'd114: q = 32'hee96d2b4;
	8'd115: q = 32'h9b919e1b;
	8'd116: q = 32'hc0c54f80;
	8'd117: q = 32'hdc20a261;
	8'd118: q = 32'h774b695a;
	8'd119: q = 32'h121a161c;
	8'd120: q = 32'h93ba0ae2;
	8'd121: q = 32'ha02ae5c0;
	8'd122: q = 32'h22e0433c;
	8'd123: q = 32'h1b171d12;
	8'd124: q = 32'h90d0b0e;
	8'd125: q = 32'h8bc7adf2;
	8'd126: q = 32'hb6a8b92d;
	8'd127: q = 32'h1ea9c814;
	8'd128: q = 32'hf1198557;
	8'd129: q = 32'h75074caf;
	8'd130: q = 32'h99ddbbee;
	8'd131: q = 32'h7f60fda3;
	8'd132: q = 32'h1269ff7;
	8'd133: q = 32'h72f5bc5c;
	8'd134: q = 32'h663bc544;
	8'd135: q = 32'hfb7e345b;
	8'd136: q = 32'h4329768b;
	8'd137: q = 32'h23c6dccb;
	8'd138: q = 32'hedfc68b6;
	8'd139: q = 32'he4f163b8;
	8'd140: q = 32'h31dccad7;
	8'd141: q = 32'h63851042;
	8'd142: q = 32'h97224013;
	8'd143: q = 32'hc6112084;
	8'd144: q = 32'h4a247d85;
	8'd145: q = 32'hbb3df8d2;
	8'd146: q = 32'hf93211ae;
	8'd147: q = 32'h29a16dc7;
	8'd148: q = 32'h9e2f4b1d;
	8'd149: q = 32'hb230f3dc;
	8'd150: q = 32'h8652ec0d;
	8'd151: q = 32'hc1e3d077;
	8'd152: q = 32'hb3166c2b;
	8'd153: q = 32'h70b999a9;
	8'd154: q = 32'h9448fa11;
	8'd155: q = 32'he9642247;
	8'd156: q = 32'hfc8cc4a8;
	8'd157: q = 32'hf03f1aa0;
	8'd158: q = 32'h7d2cd856;
	8'd159: q = 32'h3390ef22;
	8'd160: q = 32'h494ec787;
	8'd161: q = 32'h38d1c1d9;
	8'd162: q = 32'hcaa2fe8c;
	8'd163: q = 32'hd40b3698;
	8'd164: q = 32'hf581cfa6;
	8'd165: q = 32'h7ade28a5;
	8'd166: q = 32'hb78e26da;
	8'd167: q = 32'hadbfa43f;
	8'd168: q = 32'h3a9de42c;
	8'd169: q = 32'h78920d50;
	8'd170: q = 32'h5fcc9b6a;
	8'd171: q = 32'h7e466254;
	8'd172: q = 32'h8d13c2f6;
	8'd173: q = 32'hd8b8e890;
	8'd174: q = 32'h39f75e2e;
	8'd175: q = 32'hc3aff582;
	8'd176: q = 32'h5d80be9f;
	8'd177: q = 32'hd0937c69;
	8'd178: q = 32'hd52da96f;
	8'd179: q = 32'h2512b3cf;
	8'd180: q = 32'hac993bc8;
	8'd181: q = 32'h187da710;
	8'd182: q = 32'h9c636ee8;
	8'd183: q = 32'h3bbb7bdb;
	8'd184: q = 32'h267809cd;
	8'd185: q = 32'h5918f46e;
	8'd186: q = 32'h9ab701ec;
	8'd187: q = 32'h4f9aa883;
	8'd188: q = 32'h956e65e6;
	8'd189: q = 32'hffe67eaa;
	8'd190: q = 32'hbccf0821;
	8'd191: q = 32'h15e8e6ef;
	8'd192: q = 32'he79bd9ba;
	8'd193: q = 32'h6f36ce4a;
	8'd194: q = 32'h9f09d4ea;
	8'd195: q = 32'hb07cd629;
	8'd196: q = 32'ha4b2af31;
	8'd197: q = 32'h3f23312a;
	8'd198: q = 32'ha59430c6;
	8'd199: q = 32'ha266c035;
	8'd200: q = 32'h4ebc3774;
	8'd201: q = 32'h82caa6fc;
	8'd202: q = 32'h90d0b0e0;
	8'd203: q = 32'ha7d81533;
	8'd204: q = 32'h4984af1;
	8'd205: q = 32'hecdaf741;
	8'd206: q = 32'hcd500e7f;
	8'd207: q = 32'h91f62f17;
	8'd208: q = 32'h4dd68d76;
	8'd209: q = 32'hefb04d43;
	8'd210: q = 32'haa4d54cc;
	8'd211: q = 32'h9604dfe4;
	8'd212: q = 32'hd1b5e39e;
	8'd213: q = 32'h6a881b4c;
	8'd214: q = 32'h2c1fb8c1;
	8'd215: q = 32'h65517f46;
	8'd216: q = 32'h5eea049d;
	8'd217: q = 32'h8c355d01;
	8'd218: q = 32'h877473fa;
	8'd219: q = 32'hb412efb;
	8'd220: q = 32'h671d5ab3;
	8'd221: q = 32'hdbd25292;
	8'd222: q = 32'h105633e9;
	8'd223: q = 32'hd647136d;
	8'd224: q = 32'hd7618c9a;
	8'd225: q = 32'ha10c7a37;
	8'd226: q = 32'hf8148e59;
	8'd227: q = 32'h133c89eb;
	8'd228: q = 32'ha927eece;
	8'd229: q = 32'h61c935b7;
	8'd230: q = 32'h1ce5ede1;
	8'd231: q = 32'h47b13c7a;
	8'd232: q = 32'hd2df599c;
	8'd233: q = 32'hf2733f55;
	8'd234: q = 32'h14ce7918;
	8'd235: q = 32'hc737bf73;
	8'd236: q = 32'hf7cdea53;
	8'd237: q = 32'hfdaa5b5f;
	8'd238: q = 32'h3d6f14df;
	8'd239: q = 32'h44db8678;
	8'd240: q = 32'haff381ca;
	8'd241: q = 32'h68c43eb9;
	8'd242: q = 32'h24342c38;
	8'd243: q = 32'ha3405fc2;
	8'd244: q = 32'h1dc37216;
	8'd245: q = 32'he2250cbc;
	8'd246: q = 32'h3c498b28;
	8'd247: q = 32'hd9541ff;
	8'd248: q = 32'ha8017139;
	8'd249: q = 32'hcb3de08;
	8'd250: q = 32'hb4e49cd8;
	8'd251: q = 32'h56c19064;
	8'd252: q = 32'hcb84617b;
	8'd253: q = 32'h32b670d5;
	8'd254: q = 32'h6c5c7448;
	8'd255: q = 32'hb85742d0;

     endcase // case (a)
endmodule

