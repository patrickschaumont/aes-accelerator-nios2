module tboxe2(input wire clk,
              input wire [7:0] a,
              output reg [31:0] q);

   always @(posedge clk)
     case (a)
	8'd0: q = 32'h63a5c663;
	8'd1: q = 32'h7c84f87c;
	8'd2: q = 32'h7799ee77;
	8'd3: q = 32'h7b8df67b;
	8'd4: q = 32'hf20dfff2;
	8'd5: q = 32'h6bbdd66b;
	8'd6: q = 32'h6fb1de6f;
	8'd7: q = 32'hc55491c5;
	8'd8: q = 32'h30506030;
	8'd9: q = 32'h1030201;
	8'd10: q = 32'h67a9ce67;
	8'd11: q = 32'h2b7d562b;
	8'd12: q = 32'hfe19e7fe;
	8'd13: q = 32'hd762b5d7;
	8'd14: q = 32'habe64dab;
	8'd15: q = 32'h769aec76;
	8'd16: q = 32'hca458fca;
	8'd17: q = 32'h829d1f82;
	8'd18: q = 32'hc94089c9;
	8'd19: q = 32'h7d87fa7d;
	8'd20: q = 32'hfa15effa;
	8'd21: q = 32'h59ebb259;
	8'd22: q = 32'h47c98e47;
	8'd23: q = 32'hf00bfbf0;
	8'd24: q = 32'hadec41ad;
	8'd25: q = 32'hd467b3d4;
	8'd26: q = 32'ha2fd5fa2;
	8'd27: q = 32'hafea45af;
	8'd28: q = 32'h9cbf239c;
	8'd29: q = 32'ha4f753a4;
	8'd30: q = 32'h7296e472;
	8'd31: q = 32'hc05b9bc0;
	8'd32: q = 32'hb7c275b7;
	8'd33: q = 32'hfd1ce1fd;
	8'd34: q = 32'h93ae3d93;
	8'd35: q = 32'h266a4c26;
	8'd36: q = 32'h365a6c36;
	8'd37: q = 32'h3f417e3f;
	8'd38: q = 32'hf702f5f7;
	8'd39: q = 32'hcc4f83cc;
	8'd40: q = 32'h345c6834;
	8'd41: q = 32'ha5f451a5;
	8'd42: q = 32'he534d1e5;
	8'd43: q = 32'hf108f9f1;
	8'd44: q = 32'h7193e271;
	8'd45: q = 32'hd873abd8;
	8'd46: q = 32'h31536231;
	8'd47: q = 32'h153f2a15;
	8'd48: q = 32'h40c0804;
	8'd49: q = 32'hc75295c7;
	8'd50: q = 32'h23654623;
	8'd51: q = 32'hc35e9dc3;
	8'd52: q = 32'h18283018;
	8'd53: q = 32'h96a13796;
	8'd54: q = 32'h50f0a05;
	8'd55: q = 32'h9ab52f9a;
	8'd56: q = 32'h7090e07;
	8'd57: q = 32'h12362412;
	8'd58: q = 32'h809b1b80;
	8'd59: q = 32'he23ddfe2;
	8'd60: q = 32'heb26cdeb;
	8'd61: q = 32'h27694e27;
	8'd62: q = 32'hb2cd7fb2;
	8'd63: q = 32'h759fea75;
	8'd64: q = 32'h91b1209;
	8'd65: q = 32'h839e1d83;
	8'd66: q = 32'h2c74582c;
	8'd67: q = 32'h1a2e341a;
	8'd68: q = 32'h1b2d361b;
	8'd69: q = 32'h6eb2dc6e;
	8'd70: q = 32'h5aeeb45a;
	8'd71: q = 32'ha0fb5ba0;
	8'd72: q = 32'h52f6a452;
	8'd73: q = 32'h3b4d763b;
	8'd74: q = 32'hd661b7d6;
	8'd75: q = 32'hb3ce7db3;
	8'd76: q = 32'h297b5229;
	8'd77: q = 32'he33edde3;
	8'd78: q = 32'h2f715e2f;
	8'd79: q = 32'h84971384;
	8'd80: q = 32'h53f5a653;
	8'd81: q = 32'hd168b9d1;
	8'd82: q = 32'h0;
	8'd83: q = 32'hed2cc1ed;
	8'd84: q = 32'h20604020;
	8'd85: q = 32'hfc1fe3fc;
	8'd86: q = 32'hb1c879b1;
	8'd87: q = 32'h5bedb65b;
	8'd88: q = 32'h6abed46a;
	8'd89: q = 32'hcb468dcb;
	8'd90: q = 32'hbed967be;
	8'd91: q = 32'h394b7239;
	8'd92: q = 32'h4ade944a;
	8'd93: q = 32'h4cd4984c;
	8'd94: q = 32'h58e8b058;
	8'd95: q = 32'hcf4a85cf;
	8'd96: q = 32'hd06bbbd0;
	8'd97: q = 32'hef2ac5ef;
	8'd98: q = 32'haae54faa;
	8'd99: q = 32'hfb16edfb;
	8'd100: q = 32'h43c58643;
	8'd101: q = 32'h4dd79a4d;
	8'd102: q = 32'h33556633;
	8'd103: q = 32'h85941185;
	8'd104: q = 32'h45cf8a45;
	8'd105: q = 32'hf910e9f9;
	8'd106: q = 32'h2060402;
	8'd107: q = 32'h7f81fe7f;
	8'd108: q = 32'h50f0a050;
	8'd109: q = 32'h3c44783c;
	8'd110: q = 32'h9fba259f;
	8'd111: q = 32'ha8e34ba8;
	8'd112: q = 32'h51f3a251;
	8'd113: q = 32'ha3fe5da3;
	8'd114: q = 32'h40c08040;
	8'd115: q = 32'h8f8a058f;
	8'd116: q = 32'h92ad3f92;
	8'd117: q = 32'h9dbc219d;
	8'd118: q = 32'h38487038;
	8'd119: q = 32'hf504f1f5;
	8'd120: q = 32'hbcdf63bc;
	8'd121: q = 32'hb6c177b6;
	8'd122: q = 32'hda75afda;
	8'd123: q = 32'h21634221;
	8'd124: q = 32'h10302010;
	8'd125: q = 32'hff1ae5ff;
	8'd126: q = 32'hf30efdf3;
	8'd127: q = 32'hd26dbfd2;
	8'd128: q = 32'hcd4c81cd;
	8'd129: q = 32'hc14180c;
	8'd130: q = 32'h13352613;
	8'd131: q = 32'hec2fc3ec;
	8'd132: q = 32'h5fe1be5f;
	8'd133: q = 32'h97a23597;
	8'd134: q = 32'h44cc8844;
	8'd135: q = 32'h17392e17;
	8'd136: q = 32'hc45793c4;
	8'd137: q = 32'ha7f255a7;
	8'd138: q = 32'h7e82fc7e;
	8'd139: q = 32'h3d477a3d;
	8'd140: q = 32'h64acc864;
	8'd141: q = 32'h5de7ba5d;
	8'd142: q = 32'h192b3219;
	8'd143: q = 32'h7395e673;
	8'd144: q = 32'h60a0c060;
	8'd145: q = 32'h81981981;
	8'd146: q = 32'h4fd19e4f;
	8'd147: q = 32'hdc7fa3dc;
	8'd148: q = 32'h22664422;
	8'd149: q = 32'h2a7e542a;
	8'd150: q = 32'h90ab3b90;
	8'd151: q = 32'h88830b88;
	8'd152: q = 32'h46ca8c46;
	8'd153: q = 32'hee29c7ee;
	8'd154: q = 32'hb8d36bb8;
	8'd155: q = 32'h143c2814;
	8'd156: q = 32'hde79a7de;
	8'd157: q = 32'h5ee2bc5e;
	8'd158: q = 32'hb1d160b;
	8'd159: q = 32'hdb76addb;
	8'd160: q = 32'he03bdbe0;
	8'd161: q = 32'h32566432;
	8'd162: q = 32'h3a4e743a;
	8'd163: q = 32'ha1e140a;
	8'd164: q = 32'h49db9249;
	8'd165: q = 32'h60a0c06;
	8'd166: q = 32'h246c4824;
	8'd167: q = 32'h5ce4b85c;
	8'd168: q = 32'hc25d9fc2;
	8'd169: q = 32'hd36ebdd3;
	8'd170: q = 32'hacef43ac;
	8'd171: q = 32'h62a6c462;
	8'd172: q = 32'h91a83991;
	8'd173: q = 32'h95a43195;
	8'd174: q = 32'he437d3e4;
	8'd175: q = 32'h798bf279;
	8'd176: q = 32'he732d5e7;
	8'd177: q = 32'hc8438bc8;
	8'd178: q = 32'h37596e37;
	8'd179: q = 32'h6db7da6d;
	8'd180: q = 32'h8d8c018d;
	8'd181: q = 32'hd564b1d5;
	8'd182: q = 32'h4ed29c4e;
	8'd183: q = 32'ha9e049a9;
	8'd184: q = 32'h6cb4d86c;
	8'd185: q = 32'h56faac56;
	8'd186: q = 32'hf407f3f4;
	8'd187: q = 32'hea25cfea;
	8'd188: q = 32'h65afca65;
	8'd189: q = 32'h7a8ef47a;
	8'd190: q = 32'haee947ae;
	8'd191: q = 32'h8181008;
	8'd192: q = 32'hbad56fba;
	8'd193: q = 32'h7888f078;
	8'd194: q = 32'h256f4a25;
	8'd195: q = 32'h2e725c2e;
	8'd196: q = 32'h1c24381c;
	8'd197: q = 32'ha6f157a6;
	8'd198: q = 32'hb4c773b4;
	8'd199: q = 32'hc65197c6;
	8'd200: q = 32'he823cbe8;
	8'd201: q = 32'hdd7ca1dd;
	8'd202: q = 32'h749ce874;
	8'd203: q = 32'h1f213e1f;
	8'd204: q = 32'h4bdd964b;
	8'd205: q = 32'hbddc61bd;
	8'd206: q = 32'h8b860d8b;
	8'd207: q = 32'h8a850f8a;
	8'd208: q = 32'h7090e070;
	8'd209: q = 32'h3e427c3e;
	8'd210: q = 32'hb5c471b5;
	8'd211: q = 32'h66aacc66;
	8'd212: q = 32'h48d89048;
	8'd213: q = 32'h3050603;
	8'd214: q = 32'hf601f7f6;
	8'd215: q = 32'he121c0e;
	8'd216: q = 32'h61a3c261;
	8'd217: q = 32'h355f6a35;
	8'd218: q = 32'h57f9ae57;
	8'd219: q = 32'hb9d069b9;
	8'd220: q = 32'h86911786;
	8'd221: q = 32'hc15899c1;
	8'd222: q = 32'h1d273a1d;
	8'd223: q = 32'h9eb9279e;
	8'd224: q = 32'he138d9e1;
	8'd225: q = 32'hf813ebf8;
	8'd226: q = 32'h98b32b98;
	8'd227: q = 32'h11332211;
	8'd228: q = 32'h69bbd269;
	8'd229: q = 32'hd970a9d9;
	8'd230: q = 32'h8e89078e;
	8'd231: q = 32'h94a73394;
	8'd232: q = 32'h9bb62d9b;
	8'd233: q = 32'h1e223c1e;
	8'd234: q = 32'h87921587;
	8'd235: q = 32'he920c9e9;
	8'd236: q = 32'hce4987ce;
	8'd237: q = 32'h55ffaa55;
	8'd238: q = 32'h28785028;
	8'd239: q = 32'hdf7aa5df;
	8'd240: q = 32'h8c8f038c;
	8'd241: q = 32'ha1f859a1;
	8'd242: q = 32'h89800989;
	8'd243: q = 32'hd171a0d;
	8'd244: q = 32'hbfda65bf;
	8'd245: q = 32'he631d7e6;
	8'd246: q = 32'h42c68442;
	8'd247: q = 32'h68b8d068;
	8'd248: q = 32'h41c38241;
	8'd249: q = 32'h99b02999;
	8'd250: q = 32'h2d775a2d;
	8'd251: q = 32'hf111e0f;
	8'd252: q = 32'hb0cb7bb0;
	8'd253: q = 32'h54fca854;
	8'd254: q = 32'hbbd66dbb;
	8'd255: q = 32'h163a2c16;

     endcase // case (a)
endmodule

