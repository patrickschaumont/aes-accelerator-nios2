module tboxd0(input wire clk,
              input wire [7:0] a,
              output reg [31:0] q);

   always @(posedge clk)
     case (a)
	8'd0: q = 32'h51f4a750;
	8'd1: q = 32'h7e416553;
	8'd2: q = 32'h1a17a4c3;
	8'd3: q = 32'h3a275e96;
	8'd4: q = 32'h3bab6bcb;
	8'd5: q = 32'h1f9d45f1;
	8'd6: q = 32'hacfa58ab;
	8'd7: q = 32'h4be30393;
	8'd8: q = 32'h2030fa55;
	8'd9: q = 32'had766df6;
	8'd10: q = 32'h88cc7691;
	8'd11: q = 32'hf5024c25;
	8'd12: q = 32'h4fe5d7fc;
	8'd13: q = 32'hc52acbd7;
	8'd14: q = 32'h26354480;
	8'd15: q = 32'hb562a38f;
	8'd16: q = 32'hdeb15a49;
	8'd17: q = 32'h25ba1b67;
	8'd18: q = 32'h45ea0e98;
	8'd19: q = 32'h5dfec0e1;
	8'd20: q = 32'hc32f7502;
	8'd21: q = 32'h814cf012;
	8'd22: q = 32'h8d4697a3;
	8'd23: q = 32'h6bd3f9c6;
	8'd24: q = 32'h38f5fe7;
	8'd25: q = 32'h15929c95;
	8'd26: q = 32'hbf6d7aeb;
	8'd27: q = 32'h955259da;
	8'd28: q = 32'hd4be832d;
	8'd29: q = 32'h587421d3;
	8'd30: q = 32'h49e06929;
	8'd31: q = 32'h8ec9c844;
	8'd32: q = 32'h75c2896a;
	8'd33: q = 32'hf48e7978;
	8'd34: q = 32'h99583e6b;
	8'd35: q = 32'h27b971dd;
	8'd36: q = 32'hbee14fb6;
	8'd37: q = 32'hf088ad17;
	8'd38: q = 32'hc920ac66;
	8'd39: q = 32'h7dce3ab4;
	8'd40: q = 32'h63df4a18;
	8'd41: q = 32'he51a3182;
	8'd42: q = 32'h97513360;
	8'd43: q = 32'h62537f45;
	8'd44: q = 32'hb16477e0;
	8'd45: q = 32'hbb6bae84;
	8'd46: q = 32'hfe81a01c;
	8'd47: q = 32'hf9082b94;
	8'd48: q = 32'h70486858;
	8'd49: q = 32'h8f45fd19;
	8'd50: q = 32'h94de6c87;
	8'd51: q = 32'h527bf8b7;
	8'd52: q = 32'hab73d323;
	8'd53: q = 32'h724b02e2;
	8'd54: q = 32'he31f8f57;
	8'd55: q = 32'h6655ab2a;
	8'd56: q = 32'hb2eb2807;
	8'd57: q = 32'h2fb5c203;
	8'd58: q = 32'h86c57b9a;
	8'd59: q = 32'hd33708a5;
	8'd60: q = 32'h302887f2;
	8'd61: q = 32'h23bfa5b2;
	8'd62: q = 32'h2036aba;
	8'd63: q = 32'hed16825c;
	8'd64: q = 32'h8acf1c2b;
	8'd65: q = 32'ha779b492;
	8'd66: q = 32'hf307f2f0;
	8'd67: q = 32'h4e69e2a1;
	8'd68: q = 32'h65daf4cd;
	8'd69: q = 32'h605bed5;
	8'd70: q = 32'hd134621f;
	8'd71: q = 32'hc4a6fe8a;
	8'd72: q = 32'h342e539d;
	8'd73: q = 32'ha2f355a0;
	8'd74: q = 32'h58ae132;
	8'd75: q = 32'ha4f6eb75;
	8'd76: q = 32'hb83ec39;
	8'd77: q = 32'h4060efaa;
	8'd78: q = 32'h5e719f06;
	8'd79: q = 32'hbd6e1051;
	8'd80: q = 32'h3e218af9;
	8'd81: q = 32'h96dd063d;
	8'd82: q = 32'hdd3e05ae;
	8'd83: q = 32'h4de6bd46;
	8'd84: q = 32'h91548db5;
	8'd85: q = 32'h71c45d05;
	8'd86: q = 32'h406d46f;
	8'd87: q = 32'h605015ff;
	8'd88: q = 32'h1998fb24;
	8'd89: q = 32'hd6bde997;
	8'd90: q = 32'h894043cc;
	8'd91: q = 32'h67d99e77;
	8'd92: q = 32'hb0e842bd;
	8'd93: q = 32'h7898b88;
	8'd94: q = 32'he7195b38;
	8'd95: q = 32'h79c8eedb;
	8'd96: q = 32'ha17c0a47;
	8'd97: q = 32'h7c420fe9;
	8'd98: q = 32'hf8841ec9;
	8'd99: q = 32'h0;
	8'd100: q = 32'h9808683;
	8'd101: q = 32'h322bed48;
	8'd102: q = 32'h1e1170ac;
	8'd103: q = 32'h6c5a724e;
	8'd104: q = 32'hfd0efffb;
	8'd105: q = 32'hf853856;
	8'd106: q = 32'h3daed51e;
	8'd107: q = 32'h362d3927;
	8'd108: q = 32'ha0fd964;
	8'd109: q = 32'h685ca621;
	8'd110: q = 32'h9b5b54d1;
	8'd111: q = 32'h24362e3a;
	8'd112: q = 32'hc0a67b1;
	8'd113: q = 32'h9357e70f;
	8'd114: q = 32'hb4ee96d2;
	8'd115: q = 32'h1b9b919e;
	8'd116: q = 32'h80c0c54f;
	8'd117: q = 32'h61dc20a2;
	8'd118: q = 32'h5a774b69;
	8'd119: q = 32'h1c121a16;
	8'd120: q = 32'he293ba0a;
	8'd121: q = 32'hc0a02ae5;
	8'd122: q = 32'h3c22e043;
	8'd123: q = 32'h121b171d;
	8'd124: q = 32'he090d0b;
	8'd125: q = 32'hf28bc7ad;
	8'd126: q = 32'h2db6a8b9;
	8'd127: q = 32'h141ea9c8;
	8'd128: q = 32'h57f11985;
	8'd129: q = 32'haf75074c;
	8'd130: q = 32'hee99ddbb;
	8'd131: q = 32'ha37f60fd;
	8'd132: q = 32'hf701269f;
	8'd133: q = 32'h5c72f5bc;
	8'd134: q = 32'h44663bc5;
	8'd135: q = 32'h5bfb7e34;
	8'd136: q = 32'h8b432976;
	8'd137: q = 32'hcb23c6dc;
	8'd138: q = 32'hb6edfc68;
	8'd139: q = 32'hb8e4f163;
	8'd140: q = 32'hd731dcca;
	8'd141: q = 32'h42638510;
	8'd142: q = 32'h13972240;
	8'd143: q = 32'h84c61120;
	8'd144: q = 32'h854a247d;
	8'd145: q = 32'hd2bb3df8;
	8'd146: q = 32'haef93211;
	8'd147: q = 32'hc729a16d;
	8'd148: q = 32'h1d9e2f4b;
	8'd149: q = 32'hdcb230f3;
	8'd150: q = 32'hd8652ec;
	8'd151: q = 32'h77c1e3d0;
	8'd152: q = 32'h2bb3166c;
	8'd153: q = 32'ha970b999;
	8'd154: q = 32'h119448fa;
	8'd155: q = 32'h47e96422;
	8'd156: q = 32'ha8fc8cc4;
	8'd157: q = 32'ha0f03f1a;
	8'd158: q = 32'h567d2cd8;
	8'd159: q = 32'h223390ef;
	8'd160: q = 32'h87494ec7;
	8'd161: q = 32'hd938d1c1;
	8'd162: q = 32'h8ccaa2fe;
	8'd163: q = 32'h98d40b36;
	8'd164: q = 32'ha6f581cf;
	8'd165: q = 32'ha57ade28;
	8'd166: q = 32'hdab78e26;
	8'd167: q = 32'h3fadbfa4;
	8'd168: q = 32'h2c3a9de4;
	8'd169: q = 32'h5078920d;
	8'd170: q = 32'h6a5fcc9b;
	8'd171: q = 32'h547e4662;
	8'd172: q = 32'hf68d13c2;
	8'd173: q = 32'h90d8b8e8;
	8'd174: q = 32'h2e39f75e;
	8'd175: q = 32'h82c3aff5;
	8'd176: q = 32'h9f5d80be;
	8'd177: q = 32'h69d0937c;
	8'd178: q = 32'h6fd52da9;
	8'd179: q = 32'hcf2512b3;
	8'd180: q = 32'hc8ac993b;
	8'd181: q = 32'h10187da7;
	8'd182: q = 32'he89c636e;
	8'd183: q = 32'hdb3bbb7b;
	8'd184: q = 32'hcd267809;
	8'd185: q = 32'h6e5918f4;
	8'd186: q = 32'hec9ab701;
	8'd187: q = 32'h834f9aa8;
	8'd188: q = 32'he6956e65;
	8'd189: q = 32'haaffe67e;
	8'd190: q = 32'h21bccf08;
	8'd191: q = 32'hef15e8e6;
	8'd192: q = 32'hbae79bd9;
	8'd193: q = 32'h4a6f36ce;
	8'd194: q = 32'hea9f09d4;
	8'd195: q = 32'h29b07cd6;
	8'd196: q = 32'h31a4b2af;
	8'd197: q = 32'h2a3f2331;
	8'd198: q = 32'hc6a59430;
	8'd199: q = 32'h35a266c0;
	8'd200: q = 32'h744ebc37;
	8'd201: q = 32'hfc82caa6;
	8'd202: q = 32'he090d0b0;
	8'd203: q = 32'h33a7d815;
	8'd204: q = 32'hf104984a;
	8'd205: q = 32'h41ecdaf7;
	8'd206: q = 32'h7fcd500e;
	8'd207: q = 32'h1791f62f;
	8'd208: q = 32'h764dd68d;
	8'd209: q = 32'h43efb04d;
	8'd210: q = 32'hccaa4d54;
	8'd211: q = 32'he49604df;
	8'd212: q = 32'h9ed1b5e3;
	8'd213: q = 32'h4c6a881b;
	8'd214: q = 32'hc12c1fb8;
	8'd215: q = 32'h4665517f;
	8'd216: q = 32'h9d5eea04;
	8'd217: q = 32'h18c355d;
	8'd218: q = 32'hfa877473;
	8'd219: q = 32'hfb0b412e;
	8'd220: q = 32'hb3671d5a;
	8'd221: q = 32'h92dbd252;
	8'd222: q = 32'he9105633;
	8'd223: q = 32'h6dd64713;
	8'd224: q = 32'h9ad7618c;
	8'd225: q = 32'h37a10c7a;
	8'd226: q = 32'h59f8148e;
	8'd227: q = 32'heb133c89;
	8'd228: q = 32'hcea927ee;
	8'd229: q = 32'hb761c935;
	8'd230: q = 32'he11ce5ed;
	8'd231: q = 32'h7a47b13c;
	8'd232: q = 32'h9cd2df59;
	8'd233: q = 32'h55f2733f;
	8'd234: q = 32'h1814ce79;
	8'd235: q = 32'h73c737bf;
	8'd236: q = 32'h53f7cdea;
	8'd237: q = 32'h5ffdaa5b;
	8'd238: q = 32'hdf3d6f14;
	8'd239: q = 32'h7844db86;
	8'd240: q = 32'hcaaff381;
	8'd241: q = 32'hb968c43e;
	8'd242: q = 32'h3824342c;
	8'd243: q = 32'hc2a3405f;
	8'd244: q = 32'h161dc372;
	8'd245: q = 32'hbce2250c;
	8'd246: q = 32'h283c498b;
	8'd247: q = 32'hff0d9541;
	8'd248: q = 32'h39a80171;
	8'd249: q = 32'h80cb3de;
	8'd250: q = 32'hd8b4e49c;
	8'd251: q = 32'h6456c190;
	8'd252: q = 32'h7bcb8461;
	8'd253: q = 32'hd532b670;
	8'd254: q = 32'h486c5c74;
	8'd255: q = 32'hd0b85742;

     endcase // case (a)
endmodule

