
module softcore_top (
	clk_clk,
	reset_reset_n,
	pio_export);	

	input		clk_clk;
	input		reset_reset_n;
	output	[7:0]	pio_export;
endmodule
